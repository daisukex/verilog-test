module test (
  input aaa,
  input bbb,
  output ccc
);

assign ccc = aaa & bbb;

endmodule
